`ifndef INTERFACE
`define INTERFACE
//compiler directive

interface intf();
endinterface

`endif
