`ifndef DUT_TOP
`define DUT_TOP

`include "alu_simple_bugs_enc2.svp"

`endif
